module xor (input a, b, output y)
  
